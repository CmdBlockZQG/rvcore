module MUL_wallace #(XLEN = 32) (
  input clock, reset,

  input flush,

  output in_ready,
  input in_valid,
  input [1:0] in_sign,
  input [XLEN-1:0] in_a, in_b,

  input out_ready,
  output out_valid,
  output [XLEN*2-1:0] out_prod
);

  parameter YLEN = XLEN + 2; // 拓展两个符号位的位宽

  wire [YLEN-1:0] a = {{2{in_sign[1] & in_a[XLEN-1]}}, in_a};
  wire [YLEN-1:0] b = {{2{in_sign[0] & in_b[XLEN-1]}}, in_b};

  // -------------------- 部分积生成 --------------------

  reg [YLEN+1:0] p [1:YLEN/2-1];
  reg [1:0] c [YLEN/2-1]; // 最后一个部分积的减法修正必然是0

  reg [YLEN+3:0] p0;
  always_comb begin
    case (b[1:0])
      2'b00: begin // 0
        p0 = {1'b1, {YLEN+3{1'b0}}};
        c[0] = 2'b00;
      end
      2'b01: begin // +1
        p0 = {~a[YLEN-1], {3{a[YLEN-1]}}, a};
        c[0] = 2'b00;
      end
      2'b10: begin // -2
        p0 = {a[YLEN-1], {2{~a[YLEN-1]}}, ~a, 1'b0};
        c[0] = 2'b10;
      end
      2'b11: begin // -1
        p0 = {a[YLEN-1], {3{~a[YLEN-1]}}, ~a};
        c[0] = 2'b01;
      end
      default: ;
    endcase
  end

  generate
    genvar i;
    for (i = 2; i < YLEN; i = i + 2) begin : g_pi
      always_comb begin
        case (b[i+1:i-1])
          3'b000, 3'b111: begin // 0
            p[i/2] = {1'b1, {YLEN+1{1'b0}}};
            if (i != YLEN-2) c[i/2] = 2'b00;
          end
          3'b001, 3'b010: begin // +1
            p[i/2] = {~a[YLEN-1], a[YLEN-1], a};
            if (i != YLEN-2) c[i/2] = 2'b00;
          end
          3'b011: begin // +2
            p[i/2] = {~a[YLEN-1], a, 1'b0};
            if (i != YLEN-2) c[i/2] = 2'b00;
          end
          3'b100: begin // -2
            p[i/2] = {a[YLEN-1], ~a, 1'b0};
            if (i != YLEN-2) c[i/2] = 2'b10;
          end
          3'b101, 3'b110: begin // -1
            p[i/2] = {a[YLEN-1], ~a[YLEN-1], ~a};
            if (i != YLEN-2) c[i/2] = 2'b01;
          end
          default: ;
        endcase
      end
    end
  endgenerate

  // -------------------- 部分积加和测试 --------------------
  /*
  wire [2*YLEN-1:0] prod_sum [YLEN/2];
  generate
    genvar j;
    assign prod_sum[0] = {{YLEN-4{1'b0}}, p0};
    for (j = 1; j < YLEN/2; j = j + 1) begin : g_sum
      if (j == YLEN/2-1) begin : g_sum_l
        assign prod_sum[j] = {p[j], c[j-1], {((j-1)*2){1'b0}}};
      end else begin : g_sum_i
        assign prod_sum[j] = {{YLEN-3-2*j{1'b0}}, 1'b1, p[j], c[j-1], {((j-1)*2){1'b0}}};
      end
    end
  endgenerate

  reg [2*YLEN-1:0] prod;
  integer k;
  always_comb begin
    prod = 0;
    for (k = 0; k < YLEN/2; k = k + 1) begin
      prod = prod + prod_sum[k];
    end
  end
  */
  // -------------------- 华莱士树 --------------------

  ha ha_0 (.a(c[0][0]), .b(p0[0]), .s(w[0]), .cout(w[1]));
  fa fa_0 (.a(w[1]), .b(c[0][1]), .cin(p0[1]), .s(w[2]), .cout(w[3]));
  fa fa_1 (.a(w[3]), .b(c[1][0]), .cin(p[1][0]), .s(w[4]), .cout(w[5]));
  fa fa_2 (.a(w[5]), .b(c[1][1]), .cin(p[1][1]), .s(w[6]), .cout(w[7]));
  fa fa_3 (.a(w[7]), .b(c[2][0]), .cin(p[2][0]), .s(w[8]), .cout(w[9]));
  ha ha_1 (.a(p[1][2]), .b(p0[4]), .s(w[10]), .cout(w[11]));
  fa fa_4 (.a(w[11]), .b(w[9]), .cin(c[2][1]), .s(w[12]), .cout(w[13]));
  fa fa_5 (.a(p[2][1]), .b(p[1][3]), .cin(p0[5]), .s(w[14]), .cout(w[15]));
  fa fa_6 (.a(w[15]), .b(w[13]), .cin(c[3][0]), .s(w[16]), .cout(w[17]));
  fa fa_7 (.a(p[3][0]), .b(p[2][2]), .cin(p[1][4]), .s(w[18]), .cout(w[19]));
  fa fa_8 (.a(w[19]), .b(w[17]), .cin(c[3][1]), .s(w[20]), .cout(w[21]));
  fa fa_9 (.a(p[3][1]), .b(p[2][3]), .cin(p[1][5]), .s(w[22]), .cout(w[23]));
  fa fa_10 (.a(w[23]), .b(w[21]), .cin(c[4][0]), .s(w[24]), .cout(w[25]));
  fa fa_11 (.a(p[4][0]), .b(p[3][2]), .cin(p[2][4]), .s(w[26]), .cout(w[27]));
  ha ha_2 (.a(p[1][6]), .b(p0[8]), .s(w[28]), .cout(w[29]));
  fa fa_12 (.a(w[29]), .b(w[27]), .cin(w[25]), .s(w[30]), .cout(w[31]));
  fa fa_13 (.a(c[4][1]), .b(p[4][1]), .cin(p[3][3]), .s(w[32]), .cout(w[33]));
  fa fa_14 (.a(p[2][5]), .b(p[1][7]), .cin(p0[9]), .s(w[34]), .cout(w[35]));
  fa fa_15 (.a(w[35]), .b(w[33]), .cin(w[31]), .s(w[36]), .cout(w[37]));
  fa fa_16 (.a(c[5][0]), .b(p[5][0]), .cin(p[4][2]), .s(w[38]), .cout(w[39]));
  fa fa_17 (.a(p[3][4]), .b(p[2][6]), .cin(p[1][8]), .s(w[40]), .cout(w[41]));
  fa fa_18 (.a(w[41]), .b(w[39]), .cin(w[37]), .s(w[42]), .cout(w[43]));
  fa fa_19 (.a(c[5][1]), .b(p[5][1]), .cin(p[4][3]), .s(w[44]), .cout(w[45]));
  fa fa_20 (.a(p[3][5]), .b(p[2][7]), .cin(p[1][9]), .s(w[46]), .cout(w[47]));
  fa fa_21 (.a(w[47]), .b(w[45]), .cin(w[43]), .s(w[48]), .cout(w[49]));
  fa fa_22 (.a(c[6][0]), .b(p[6][0]), .cin(p[5][2]), .s(w[50]), .cout(w[51]));
  fa fa_23 (.a(p[4][4]), .b(p[3][6]), .cin(p[2][8]), .s(w[52]), .cout(w[53]));
  ha ha_3 (.a(p[1][10]), .b(p0[12]), .s(w[54]), .cout(w[55]));
  fa fa_24 (.a(w[55]), .b(w[53]), .cin(w[51]), .s(w[56]), .cout(w[57]));
  fa fa_25 (.a(w[49]), .b(c[6][1]), .cin(p[6][1]), .s(w[58]), .cout(w[59]));
  fa fa_26 (.a(p[5][3]), .b(p[4][5]), .cin(p[3][7]), .s(w[60]), .cout(w[61]));
  fa fa_27 (.a(p[2][9]), .b(p[1][11]), .cin(p0[13]), .s(w[62]), .cout(w[63]));
  fa fa_28 (.a(w[63]), .b(w[61]), .cin(w[59]), .s(w[64]), .cout(w[65]));
  fa fa_29 (.a(w[57]), .b(c[7][0]), .cin(p[7][0]), .s(w[66]), .cout(w[67]));
  fa fa_30 (.a(p[6][2]), .b(p[5][4]), .cin(p[4][6]), .s(w[68]), .cout(w[69]));
  fa fa_31 (.a(p[3][8]), .b(p[2][10]), .cin(p[1][12]), .s(w[70]), .cout(w[71]));
  fa fa_32 (.a(w[71]), .b(w[69]), .cin(w[67]), .s(w[72]), .cout(w[73]));
  fa fa_33 (.a(w[65]), .b(c[7][1]), .cin(p[7][1]), .s(w[74]), .cout(w[75]));
  fa fa_34 (.a(p[6][3]), .b(p[5][5]), .cin(p[4][7]), .s(w[76]), .cout(w[77]));
  fa fa_35 (.a(p[3][9]), .b(p[2][11]), .cin(p[1][13]), .s(w[78]), .cout(w[79]));
  fa fa_36 (.a(w[79]), .b(w[77]), .cin(w[75]), .s(w[80]), .cout(w[81]));
  fa fa_37 (.a(w[73]), .b(c[8][0]), .cin(p[8][0]), .s(w[82]), .cout(w[83]));
  fa fa_38 (.a(p[7][2]), .b(p[6][4]), .cin(p[5][6]), .s(w[84]), .cout(w[85]));
  fa fa_39 (.a(p[4][8]), .b(p[3][10]), .cin(p[2][12]), .s(w[86]), .cout(w[87]));
  ha ha_4 (.a(p[1][14]), .b(p0[16]), .s(w[88]), .cout(w[89]));
  fa fa_40 (.a(w[89]), .b(w[87]), .cin(w[85]), .s(w[90]), .cout(w[91]));
  fa fa_41 (.a(w[83]), .b(w[81]), .cin(c[8][1]), .s(w[92]), .cout(w[93]));
  fa fa_42 (.a(p[8][1]), .b(p[7][3]), .cin(p[6][5]), .s(w[94]), .cout(w[95]));
  fa fa_43 (.a(p[5][7]), .b(p[4][9]), .cin(p[3][11]), .s(w[96]), .cout(w[97]));
  fa fa_44 (.a(p[2][13]), .b(p[1][15]), .cin(p0[17]), .s(w[98]), .cout(w[99]));
  fa fa_45 (.a(w[99]), .b(w[97]), .cin(w[95]), .s(w[100]), .cout(w[101]));
  fa fa_46 (.a(w[93]), .b(w[91]), .cin(c[9][0]), .s(w[102]), .cout(w[103]));
  fa fa_47 (.a(p[9][0]), .b(p[8][2]), .cin(p[7][4]), .s(w[104]), .cout(w[105]));
  fa fa_48 (.a(p[6][6]), .b(p[5][8]), .cin(p[4][10]), .s(w[106]), .cout(w[107]));
  fa fa_49 (.a(p[3][12]), .b(p[2][14]), .cin(p[1][16]), .s(w[108]), .cout(w[109]));
  fa fa_50 (.a(w[109]), .b(w[107]), .cin(w[105]), .s(w[110]), .cout(w[111]));
  fa fa_51 (.a(w[103]), .b(w[101]), .cin(c[9][1]), .s(w[112]), .cout(w[113]));
  fa fa_52 (.a(p[9][1]), .b(p[8][3]), .cin(p[7][5]), .s(w[114]), .cout(w[115]));
  fa fa_53 (.a(p[6][7]), .b(p[5][9]), .cin(p[4][11]), .s(w[116]), .cout(w[117]));
  fa fa_54 (.a(p[3][13]), .b(p[2][15]), .cin(p[1][17]), .s(w[118]), .cout(w[119]));
  fa fa_55 (.a(w[119]), .b(w[117]), .cin(w[115]), .s(w[120]), .cout(w[121]));
  fa fa_56 (.a(w[113]), .b(w[111]), .cin(c[10][0]), .s(w[122]), .cout(w[123]));
  fa fa_57 (.a(p[10][0]), .b(p[9][2]), .cin(p[8][4]), .s(w[124]), .cout(w[125]));
  fa fa_58 (.a(p[7][6]), .b(p[6][8]), .cin(p[5][10]), .s(w[126]), .cout(w[127]));
  fa fa_59 (.a(p[4][12]), .b(p[3][14]), .cin(p[2][16]), .s(w[128]), .cout(w[129]));
  ha ha_5 (.a(p[1][18]), .b(p0[20]), .s(w[130]), .cout(w[131]));
  fa fa_60 (.a(w[131]), .b(w[129]), .cin(w[127]), .s(w[132]), .cout(w[133]));
  fa fa_61 (.a(w[125]), .b(w[123]), .cin(w[121]), .s(w[134]), .cout(w[135]));
  fa fa_62 (.a(c[10][1]), .b(p[10][1]), .cin(p[9][3]), .s(w[136]), .cout(w[137]));
  fa fa_63 (.a(p[8][5]), .b(p[7][7]), .cin(p[6][9]), .s(w[138]), .cout(w[139]));
  fa fa_64 (.a(p[5][11]), .b(p[4][13]), .cin(p[3][15]), .s(w[140]), .cout(w[141]));
  fa fa_65 (.a(p[2][17]), .b(p[1][19]), .cin(p0[21]), .s(w[142]), .cout(w[143]));
  fa fa_66 (.a(w[143]), .b(w[141]), .cin(w[139]), .s(w[144]), .cout(w[145]));
  fa fa_67 (.a(w[137]), .b(w[135]), .cin(w[133]), .s(w[146]), .cout(w[147]));
  fa fa_68 (.a(c[11][0]), .b(p[11][0]), .cin(p[10][2]), .s(w[148]), .cout(w[149]));
  fa fa_69 (.a(p[9][4]), .b(p[8][6]), .cin(p[7][8]), .s(w[150]), .cout(w[151]));
  fa fa_70 (.a(p[6][10]), .b(p[5][12]), .cin(p[4][14]), .s(w[152]), .cout(w[153]));
  fa fa_71 (.a(p[3][16]), .b(p[2][18]), .cin(p[1][20]), .s(w[154]), .cout(w[155]));
  fa fa_72 (.a(w[155]), .b(w[153]), .cin(w[151]), .s(w[156]), .cout(w[157]));
  fa fa_73 (.a(w[149]), .b(w[147]), .cin(w[145]), .s(w[158]), .cout(w[159]));
  fa fa_74 (.a(c[11][1]), .b(p[11][1]), .cin(p[10][3]), .s(w[160]), .cout(w[161]));
  fa fa_75 (.a(p[9][5]), .b(p[8][7]), .cin(p[7][9]), .s(w[162]), .cout(w[163]));
  fa fa_76 (.a(p[6][11]), .b(p[5][13]), .cin(p[4][15]), .s(w[164]), .cout(w[165]));
  fa fa_77 (.a(p[3][17]), .b(p[2][19]), .cin(p[1][21]), .s(w[166]), .cout(w[167]));
  fa fa_78 (.a(w[167]), .b(w[165]), .cin(w[163]), .s(w[168]), .cout(w[169]));
  fa fa_79 (.a(w[161]), .b(w[159]), .cin(w[157]), .s(w[170]), .cout(w[171]));
  fa fa_80 (.a(c[12][0]), .b(p[12][0]), .cin(p[11][2]), .s(w[172]), .cout(w[173]));
  fa fa_81 (.a(p[10][4]), .b(p[9][6]), .cin(p[8][8]), .s(w[174]), .cout(w[175]));
  fa fa_82 (.a(p[7][10]), .b(p[6][12]), .cin(p[5][14]), .s(w[176]), .cout(w[177]));
  fa fa_83 (.a(p[4][16]), .b(p[3][18]), .cin(p[2][20]), .s(w[178]), .cout(w[179]));
  ha ha_6 (.a(p[1][22]), .b(p0[24]), .s(w[180]), .cout(w[181]));
  fa fa_84 (.a(w[181]), .b(w[179]), .cin(w[177]), .s(w[182]), .cout(w[183]));
  fa fa_85 (.a(w[175]), .b(w[173]), .cin(w[171]), .s(w[184]), .cout(w[185]));
  fa fa_86 (.a(w[169]), .b(c[12][1]), .cin(p[12][1]), .s(w[186]), .cout(w[187]));
  fa fa_87 (.a(p[11][3]), .b(p[10][5]), .cin(p[9][7]), .s(w[188]), .cout(w[189]));
  fa fa_88 (.a(p[8][9]), .b(p[7][11]), .cin(p[6][13]), .s(w[190]), .cout(w[191]));
  fa fa_89 (.a(p[5][15]), .b(p[4][17]), .cin(p[3][19]), .s(w[192]), .cout(w[193]));
  fa fa_90 (.a(p[2][21]), .b(p[1][23]), .cin(p0[25]), .s(w[194]), .cout(w[195]));
  fa fa_91 (.a(w[195]), .b(w[193]), .cin(w[191]), .s(w[196]), .cout(w[197]));
  fa fa_92 (.a(w[189]), .b(w[187]), .cin(w[185]), .s(w[198]), .cout(w[199]));
  fa fa_93 (.a(w[183]), .b(c[13][0]), .cin(p[13][0]), .s(w[200]), .cout(w[201]));
  fa fa_94 (.a(p[12][2]), .b(p[11][4]), .cin(p[10][6]), .s(w[202]), .cout(w[203]));
  fa fa_95 (.a(p[9][8]), .b(p[8][10]), .cin(p[7][12]), .s(w[204]), .cout(w[205]));
  fa fa_96 (.a(p[6][14]), .b(p[5][16]), .cin(p[4][18]), .s(w[206]), .cout(w[207]));
  fa fa_97 (.a(p[3][20]), .b(p[2][22]), .cin(p[1][24]), .s(w[208]), .cout(w[209]));
  fa fa_98 (.a(w[209]), .b(w[207]), .cin(w[205]), .s(w[210]), .cout(w[211]));
  fa fa_99 (.a(w[203]), .b(w[201]), .cin(w[199]), .s(w[212]), .cout(w[213]));
  fa fa_100 (.a(w[197]), .b(c[13][1]), .cin(p[13][1]), .s(w[214]), .cout(w[215]));
  fa fa_101 (.a(p[12][3]), .b(p[11][5]), .cin(p[10][7]), .s(w[216]), .cout(w[217]));
  fa fa_102 (.a(p[9][9]), .b(p[8][11]), .cin(p[7][13]), .s(w[218]), .cout(w[219]));
  fa fa_103 (.a(p[6][15]), .b(p[5][17]), .cin(p[4][19]), .s(w[220]), .cout(w[221]));
  fa fa_104 (.a(p[3][21]), .b(p[2][23]), .cin(p[1][25]), .s(w[222]), .cout(w[223]));
  fa fa_105 (.a(w[223]), .b(w[221]), .cin(w[219]), .s(w[224]), .cout(w[225]));
  fa fa_106 (.a(w[217]), .b(w[215]), .cin(w[213]), .s(w[226]), .cout(w[227]));
  fa fa_107 (.a(w[211]), .b(c[14][0]), .cin(p[14][0]), .s(w[228]), .cout(w[229]));
  fa fa_108 (.a(p[13][2]), .b(p[12][4]), .cin(p[11][6]), .s(w[230]), .cout(w[231]));
  fa fa_109 (.a(p[10][8]), .b(p[9][10]), .cin(p[8][12]), .s(w[232]), .cout(w[233]));
  fa fa_110 (.a(p[7][14]), .b(p[6][16]), .cin(p[5][18]), .s(w[234]), .cout(w[235]));
  fa fa_111 (.a(p[4][20]), .b(p[3][22]), .cin(p[2][24]), .s(w[236]), .cout(w[237]));
  ha ha_7 (.a(p[1][26]), .b(p0[28]), .s(w[238]), .cout(w[239]));
  fa fa_112 (.a(w[239]), .b(w[237]), .cin(w[235]), .s(w[240]), .cout(w[241]));
  fa fa_113 (.a(w[233]), .b(w[231]), .cin(w[229]), .s(w[242]), .cout(w[243]));
  fa fa_114 (.a(w[227]), .b(w[225]), .cin(c[14][1]), .s(w[244]), .cout(w[245]));
  fa fa_115 (.a(p[14][1]), .b(p[13][3]), .cin(p[12][5]), .s(w[246]), .cout(w[247]));
  fa fa_116 (.a(p[11][7]), .b(p[10][9]), .cin(p[9][11]), .s(w[248]), .cout(w[249]));
  fa fa_117 (.a(p[8][13]), .b(p[7][15]), .cin(p[6][17]), .s(w[250]), .cout(w[251]));
  fa fa_118 (.a(p[5][19]), .b(p[4][21]), .cin(p[3][23]), .s(w[252]), .cout(w[253]));
  fa fa_119 (.a(p[2][25]), .b(p[1][27]), .cin(p0[29]), .s(w[254]), .cout(w[255]));
  fa fa_120 (.a(w[255]), .b(w[253]), .cin(w[251]), .s(w[256]), .cout(w[257]));
  fa fa_121 (.a(w[249]), .b(w[247]), .cin(w[245]), .s(w[258]), .cout(w[259]));
  fa fa_122 (.a(w[243]), .b(w[241]), .cin(c[15][0]), .s(w[260]), .cout(w[261]));
  fa fa_123 (.a(p[15][0]), .b(p[14][2]), .cin(p[13][4]), .s(w[262]), .cout(w[263]));
  fa fa_124 (.a(p[12][6]), .b(p[11][8]), .cin(p[10][10]), .s(w[264]), .cout(w[265]));
  fa fa_125 (.a(p[9][12]), .b(p[8][14]), .cin(p[7][16]), .s(w[266]), .cout(w[267]));
  fa fa_126 (.a(p[6][18]), .b(p[5][20]), .cin(p[4][22]), .s(w[268]), .cout(w[269]));
  fa fa_127 (.a(p[3][24]), .b(p[2][26]), .cin(p[1][28]), .s(w[270]), .cout(w[271]));
  fa fa_128 (.a(w[271]), .b(w[269]), .cin(w[267]), .s(w[272]), .cout(w[273]));
  fa fa_129 (.a(w[265]), .b(w[263]), .cin(w[261]), .s(w[274]), .cout(w[275]));
  fa fa_130 (.a(w[259]), .b(w[257]), .cin(c[15][1]), .s(w[276]), .cout(w[277]));
  fa fa_131 (.a(p[15][1]), .b(p[14][3]), .cin(p[13][5]), .s(w[278]), .cout(w[279]));
  fa fa_132 (.a(p[12][7]), .b(p[11][9]), .cin(p[10][11]), .s(w[280]), .cout(w[281]));
  fa fa_133 (.a(p[9][13]), .b(p[8][15]), .cin(p[7][17]), .s(w[282]), .cout(w[283]));
  fa fa_134 (.a(p[6][19]), .b(p[5][21]), .cin(p[4][23]), .s(w[284]), .cout(w[285]));
  fa fa_135 (.a(p[3][25]), .b(p[2][27]), .cin(p[1][29]), .s(w[286]), .cout(w[287]));
  fa fa_136 (.a(w[287]), .b(w[285]), .cin(w[283]), .s(w[288]), .cout(w[289]));
  fa fa_137 (.a(w[281]), .b(w[279]), .cin(w[277]), .s(w[290]), .cout(w[291]));
  fa fa_138 (.a(w[275]), .b(w[273]), .cin(p[16][0]), .s(w[292]), .cout(w[293]));
  fa fa_139 (.a(p[15][2]), .b(p[14][4]), .cin(p[13][6]), .s(w[294]), .cout(w[295]));
  fa fa_140 (.a(p[12][8]), .b(p[11][10]), .cin(p[10][12]), .s(w[296]), .cout(w[297]));
  fa fa_141 (.a(p[9][14]), .b(p[8][16]), .cin(p[7][18]), .s(w[298]), .cout(w[299]));
  fa fa_142 (.a(p[6][20]), .b(p[5][22]), .cin(p[4][24]), .s(w[300]), .cout(w[301]));
  fa fa_143 (.a(p[3][26]), .b(p[2][28]), .cin(p[1][30]), .s(w[302]), .cout(w[303]));
  fa fa_144 (.a(w[303]), .b(w[301]), .cin(w[299]), .s(w[304]), .cout(w[305]));
  fa fa_145 (.a(w[297]), .b(w[295]), .cin(w[293]), .s(w[306]), .cout(w[307]));
  fa fa_146 (.a(w[291]), .b(w[289]), .cin(p[16][1]), .s(w[308]), .cout(w[309]));
  fa fa_147 (.a(p[15][3]), .b(p[14][5]), .cin(p[13][7]), .s(w[310]), .cout(w[311]));
  fa fa_148 (.a(p[12][9]), .b(p[11][11]), .cin(p[10][13]), .s(w[312]), .cout(w[313]));
  fa fa_149 (.a(p[9][15]), .b(p[8][17]), .cin(p[7][19]), .s(w[314]), .cout(w[315]));
  fa fa_150 (.a(p[6][21]), .b(p[5][23]), .cin(p[4][25]), .s(w[316]), .cout(w[317]));
  fa fa_151 (.a(p[3][27]), .b(p[2][29]), .cin(p[1][31]), .s(w[318]), .cout(w[319]));
  fa fa_152 (.a(w[319]), .b(w[317]), .cin(w[315]), .s(w[320]), .cout(w[321]));
  fa fa_153 (.a(w[313]), .b(w[311]), .cin(w[309]), .s(w[322]), .cout(w[323]));
  fa fa_154 (.a(w[307]), .b(w[305]), .cin(p[16][2]), .s(w[324]), .cout(w[325]));
  fa fa_155 (.a(p[15][4]), .b(p[14][6]), .cin(p[13][8]), .s(w[326]), .cout(w[327]));
  fa fa_156 (.a(p[12][10]), .b(p[11][12]), .cin(p[10][14]), .s(w[328]), .cout(w[329]));
  fa fa_157 (.a(p[9][16]), .b(p[8][18]), .cin(p[7][20]), .s(w[330]), .cout(w[331]));
  fa fa_158 (.a(p[6][22]), .b(p[5][24]), .cin(p[4][26]), .s(w[332]), .cout(w[333]));
  fa fa_159 (.a(p[3][28]), .b(p[2][30]), .cin(p[1][32]), .s(w[334]), .cout(w[335]));
  fa fa_160 (.a(w[335]), .b(w[333]), .cin(w[331]), .s(w[336]), .cout(w[337]));
  fa fa_161 (.a(w[329]), .b(w[327]), .cin(w[325]), .s(w[338]), .cout(w[339]));
  fa fa_162 (.a(w[323]), .b(w[321]), .cin(p[16][3]), .s(w[340]), .cout(w[341]));
  fa fa_163 (.a(p[15][5]), .b(p[14][7]), .cin(p[13][9]), .s(w[342]), .cout(w[343]));
  fa fa_164 (.a(p[12][11]), .b(p[11][13]), .cin(p[10][15]), .s(w[344]), .cout(w[345]));
  fa fa_165 (.a(p[9][17]), .b(p[8][19]), .cin(p[7][21]), .s(w[346]), .cout(w[347]));
  fa fa_166 (.a(p[6][23]), .b(p[5][25]), .cin(p[4][27]), .s(w[348]), .cout(w[349]));
  fa fa_167 (.a(p[3][29]), .b(p[2][31]), .cin(p[1][33]), .s(w[350]), .cout(w[351]));
  fa fa_168 (.a(w[351]), .b(w[349]), .cin(w[347]), .s(w[352]), .cout(w[353]));
  fa fa_169 (.a(w[345]), .b(w[343]), .cin(w[341]), .s(w[354]), .cout(w[355]));
  fa fa_170 (.a(w[339]), .b(w[337]), .cin(p[16][4]), .s(w[356]), .cout(w[357]));
  fa fa_171 (.a(p[15][6]), .b(p[14][8]), .cin(p[13][10]), .s(w[358]), .cout(w[359]));
  fa fa_172 (.a(p[12][12]), .b(p[11][14]), .cin(p[10][16]), .s(w[360]), .cout(w[361]));
  fa fa_173 (.a(p[9][18]), .b(p[8][20]), .cin(p[7][22]), .s(w[362]), .cout(w[363]));
  fa fa_174 (.a(p[6][24]), .b(p[5][26]), .cin(p[4][28]), .s(w[364]), .cout(w[365]));
  fa fa_175 (.a(p[3][30]), .b(p[2][32]), .cin(p[1][34]), .s(w[366]), .cout(w[367]));
  fa fa_176 (.a(w[367]), .b(w[365]), .cin(w[363]), .s(w[368]), .cout(w[369]));
  fa fa_177 (.a(w[361]), .b(w[359]), .cin(w[357]), .s(w[370]), .cout(w[371]));
  fa fa_178 (.a(w[355]), .b(w[353]), .cin(p[16][5]), .s(w[372]), .cout(w[373]));
  fa fa_179 (.a(p[15][7]), .b(p[14][9]), .cin(p[13][11]), .s(w[374]), .cout(w[375]));
  fa fa_180 (.a(p[12][13]), .b(p[11][15]), .cin(p[10][17]), .s(w[376]), .cout(w[377]));
  fa fa_181 (.a(p[9][19]), .b(p[8][21]), .cin(p[7][23]), .s(w[378]), .cout(w[379]));
  fa fa_182 (.a(p[6][25]), .b(p[5][27]), .cin(p[4][29]), .s(w[380]), .cout(w[381]));
  fa fa_183 (.a(p[3][31]), .b(p[2][33]), .cin(p[1][35]), .s(w[382]), .cout(w[383]));
  fa fa_184 (.a(w[383]), .b(w[381]), .cin(w[379]), .s(w[384]), .cout(w[385]));
  fa fa_185 (.a(w[377]), .b(w[375]), .cin(w[373]), .s(w[386]), .cout(w[387]));
  fa fa_186 (.a(w[371]), .b(w[369]), .cin(p[16][6]), .s(w[388]), .cout(w[389]));
  fa fa_187 (.a(p[15][8]), .b(p[14][10]), .cin(p[13][12]), .s(w[390]), .cout(w[391]));
  fa fa_188 (.a(p[12][14]), .b(p[11][16]), .cin(p[10][18]), .s(w[392]), .cout(w[393]));
  fa fa_189 (.a(p[9][20]), .b(p[8][22]), .cin(p[7][24]), .s(w[394]), .cout(w[395]));
  fa fa_190 (.a(p[6][26]), .b(p[5][28]), .cin(p[4][30]), .s(w[396]), .cout(w[397]));
  fa fa_191 (.a(p[3][32]), .b(p[2][34]), .cin(1'b1), .s(w[398]), .cout(w[399]));
  fa fa_192 (.a(w[399]), .b(w[397]), .cin(w[395]), .s(w[400]), .cout(w[401]));
  fa fa_193 (.a(w[393]), .b(w[391]), .cin(w[389]), .s(w[402]), .cout(w[403]));
  fa fa_194 (.a(w[387]), .b(w[385]), .cin(p[16][7]), .s(w[404]), .cout(w[405]));
  fa fa_195 (.a(p[15][9]), .b(p[14][11]), .cin(p[13][13]), .s(w[406]), .cout(w[407]));
  fa fa_196 (.a(p[12][15]), .b(p[11][17]), .cin(p[10][19]), .s(w[408]), .cout(w[409]));
  fa fa_197 (.a(p[9][21]), .b(p[8][23]), .cin(p[7][25]), .s(w[410]), .cout(w[411]));
  fa fa_198 (.a(p[6][27]), .b(p[5][29]), .cin(p[4][31]), .s(w[412]), .cout(w[413]));
  ha ha_8 (.a(p[3][33]), .b(p[2][35]), .s(w[414]), .cout(w[415]));
  fa fa_199 (.a(w[415]), .b(w[413]), .cin(w[411]), .s(w[416]), .cout(w[417]));
  fa fa_200 (.a(w[409]), .b(w[407]), .cin(w[405]), .s(w[418]), .cout(w[419]));
  fa fa_201 (.a(w[403]), .b(w[401]), .cin(p[16][8]), .s(w[420]), .cout(w[421]));
  fa fa_202 (.a(p[15][10]), .b(p[14][12]), .cin(p[13][14]), .s(w[422]), .cout(w[423]));
  fa fa_203 (.a(p[12][16]), .b(p[11][18]), .cin(p[10][20]), .s(w[424]), .cout(w[425]));
  fa fa_204 (.a(p[9][22]), .b(p[8][24]), .cin(p[7][26]), .s(w[426]), .cout(w[427]));
  fa fa_205 (.a(p[6][28]), .b(p[5][30]), .cin(p[4][32]), .s(w[428]), .cout(w[429]));
  ha ha_9 (.a(p[3][34]), .b(1'b1), .s(w[430]), .cout(w[431]));
  fa fa_206 (.a(w[431]), .b(w[429]), .cin(w[427]), .s(w[432]), .cout(w[433]));
  fa fa_207 (.a(w[425]), .b(w[423]), .cin(w[421]), .s(w[434]), .cout(w[435]));
  fa fa_208 (.a(w[419]), .b(w[417]), .cin(p[16][9]), .s(w[436]), .cout(w[437]));
  fa fa_209 (.a(p[15][11]), .b(p[14][13]), .cin(p[13][15]), .s(w[438]), .cout(w[439]));
  fa fa_210 (.a(p[12][17]), .b(p[11][19]), .cin(p[10][21]), .s(w[440]), .cout(w[441]));
  fa fa_211 (.a(p[9][23]), .b(p[8][25]), .cin(p[7][27]), .s(w[442]), .cout(w[443]));
  fa fa_212 (.a(p[6][29]), .b(p[5][31]), .cin(p[4][33]), .s(w[444]), .cout(w[445]));
  fa fa_213 (.a(w[445]), .b(w[443]), .cin(w[441]), .s(w[446]), .cout(w[447]));
  fa fa_214 (.a(w[439]), .b(w[437]), .cin(w[435]), .s(w[448]), .cout(w[449]));
  fa fa_215 (.a(w[433]), .b(p[16][10]), .cin(p[15][12]), .s(w[450]), .cout(w[451]));
  fa fa_216 (.a(p[14][14]), .b(p[13][16]), .cin(p[12][18]), .s(w[452]), .cout(w[453]));
  fa fa_217 (.a(p[11][20]), .b(p[10][22]), .cin(p[9][24]), .s(w[454]), .cout(w[455]));
  fa fa_218 (.a(p[8][26]), .b(p[7][28]), .cin(p[6][30]), .s(w[456]), .cout(w[457]));
  fa fa_219 (.a(p[5][32]), .b(p[4][34]), .cin(1'b1), .s(w[458]), .cout(w[459]));
  fa fa_220 (.a(w[459]), .b(w[457]), .cin(w[455]), .s(w[460]), .cout(w[461]));
  fa fa_221 (.a(w[453]), .b(w[451]), .cin(w[449]), .s(w[462]), .cout(w[463]));
  fa fa_222 (.a(w[447]), .b(p[16][11]), .cin(p[15][13]), .s(w[464]), .cout(w[465]));
  fa fa_223 (.a(p[14][15]), .b(p[13][17]), .cin(p[12][19]), .s(w[466]), .cout(w[467]));
  fa fa_224 (.a(p[11][21]), .b(p[10][23]), .cin(p[9][25]), .s(w[468]), .cout(w[469]));
  fa fa_225 (.a(p[8][27]), .b(p[7][29]), .cin(p[6][31]), .s(w[470]), .cout(w[471]));
  ha ha_10 (.a(p[5][33]), .b(p[4][35]), .s(w[472]), .cout(w[473]));
  fa fa_226 (.a(w[473]), .b(w[471]), .cin(w[469]), .s(w[474]), .cout(w[475]));
  fa fa_227 (.a(w[467]), .b(w[465]), .cin(w[463]), .s(w[476]), .cout(w[477]));
  fa fa_228 (.a(w[461]), .b(p[16][12]), .cin(p[15][14]), .s(w[478]), .cout(w[479]));
  fa fa_229 (.a(p[14][16]), .b(p[13][18]), .cin(p[12][20]), .s(w[480]), .cout(w[481]));
  fa fa_230 (.a(p[11][22]), .b(p[10][24]), .cin(p[9][26]), .s(w[482]), .cout(w[483]));
  fa fa_231 (.a(p[8][28]), .b(p[7][30]), .cin(p[6][32]), .s(w[484]), .cout(w[485]));
  ha ha_11 (.a(p[5][34]), .b(1'b1), .s(w[486]), .cout(w[487]));
  fa fa_232 (.a(w[487]), .b(w[485]), .cin(w[483]), .s(w[488]), .cout(w[489]));
  fa fa_233 (.a(w[481]), .b(w[479]), .cin(w[477]), .s(w[490]), .cout(w[491]));
  fa fa_234 (.a(w[475]), .b(p[16][13]), .cin(p[15][15]), .s(w[492]), .cout(w[493]));
  fa fa_235 (.a(p[14][17]), .b(p[13][19]), .cin(p[12][21]), .s(w[494]), .cout(w[495]));
  fa fa_236 (.a(p[11][23]), .b(p[10][25]), .cin(p[9][27]), .s(w[496]), .cout(w[497]));
  fa fa_237 (.a(p[8][29]), .b(p[7][31]), .cin(p[6][33]), .s(w[498]), .cout(w[499]));
  fa fa_238 (.a(w[499]), .b(w[497]), .cin(w[495]), .s(w[500]), .cout(w[501]));
  fa fa_239 (.a(w[493]), .b(w[491]), .cin(w[489]), .s(w[502]), .cout(w[503]));
  fa fa_240 (.a(p[16][14]), .b(p[15][16]), .cin(p[14][18]), .s(w[504]), .cout(w[505]));
  fa fa_241 (.a(p[13][20]), .b(p[12][22]), .cin(p[11][24]), .s(w[506]), .cout(w[507]));
  fa fa_242 (.a(p[10][26]), .b(p[9][28]), .cin(p[8][30]), .s(w[508]), .cout(w[509]));
  fa fa_243 (.a(p[7][32]), .b(p[6][34]), .cin(1'b1), .s(w[510]), .cout(w[511]));
  fa fa_244 (.a(w[511]), .b(w[509]), .cin(w[507]), .s(w[512]), .cout(w[513]));
  fa fa_245 (.a(w[505]), .b(w[503]), .cin(w[501]), .s(w[514]), .cout(w[515]));
  fa fa_246 (.a(p[16][15]), .b(p[15][17]), .cin(p[14][19]), .s(w[516]), .cout(w[517]));
  fa fa_247 (.a(p[13][21]), .b(p[12][23]), .cin(p[11][25]), .s(w[518]), .cout(w[519]));
  fa fa_248 (.a(p[10][27]), .b(p[9][29]), .cin(p[8][31]), .s(w[520]), .cout(w[521]));
  ha ha_12 (.a(p[7][33]), .b(p[6][35]), .s(w[522]), .cout(w[523]));
  fa fa_249 (.a(w[523]), .b(w[521]), .cin(w[519]), .s(w[524]), .cout(w[525]));
  fa fa_250 (.a(w[517]), .b(w[515]), .cin(w[513]), .s(w[526]), .cout(w[527]));
  fa fa_251 (.a(p[16][16]), .b(p[15][18]), .cin(p[14][20]), .s(w[528]), .cout(w[529]));
  fa fa_252 (.a(p[13][22]), .b(p[12][24]), .cin(p[11][26]), .s(w[530]), .cout(w[531]));
  fa fa_253 (.a(p[10][28]), .b(p[9][30]), .cin(p[8][32]), .s(w[532]), .cout(w[533]));
  ha ha_13 (.a(p[7][34]), .b(1'b1), .s(w[534]), .cout(w[535]));
  fa fa_254 (.a(w[535]), .b(w[533]), .cin(w[531]), .s(w[536]), .cout(w[537]));
  fa fa_255 (.a(w[529]), .b(w[527]), .cin(w[525]), .s(w[538]), .cout(w[539]));
  fa fa_256 (.a(p[16][17]), .b(p[15][19]), .cin(p[14][21]), .s(w[540]), .cout(w[541]));
  fa fa_257 (.a(p[13][23]), .b(p[12][25]), .cin(p[11][27]), .s(w[542]), .cout(w[543]));
  fa fa_258 (.a(p[10][29]), .b(p[9][31]), .cin(p[8][33]), .s(w[544]), .cout(w[545]));
  fa fa_259 (.a(w[545]), .b(w[543]), .cin(w[541]), .s(w[546]), .cout(w[547]));
  fa fa_260 (.a(w[539]), .b(w[537]), .cin(p[16][18]), .s(w[548]), .cout(w[549]));
  fa fa_261 (.a(p[15][20]), .b(p[14][22]), .cin(p[13][24]), .s(w[550]), .cout(w[551]));
  fa fa_262 (.a(p[12][26]), .b(p[11][28]), .cin(p[10][30]), .s(w[552]), .cout(w[553]));
  fa fa_263 (.a(p[9][32]), .b(p[8][34]), .cin(1'b1), .s(w[554]), .cout(w[555]));
  fa fa_264 (.a(w[555]), .b(w[553]), .cin(w[551]), .s(w[556]), .cout(w[557]));
  fa fa_265 (.a(w[549]), .b(w[547]), .cin(p[16][19]), .s(w[558]), .cout(w[559]));
  fa fa_266 (.a(p[15][21]), .b(p[14][23]), .cin(p[13][25]), .s(w[560]), .cout(w[561]));
  fa fa_267 (.a(p[12][27]), .b(p[11][29]), .cin(p[10][31]), .s(w[562]), .cout(w[563]));
  ha ha_14 (.a(p[9][33]), .b(p[8][35]), .s(w[564]), .cout(w[565]));
  fa fa_268 (.a(w[565]), .b(w[563]), .cin(w[561]), .s(w[566]), .cout(w[567]));
  fa fa_269 (.a(w[559]), .b(w[557]), .cin(p[16][20]), .s(w[568]), .cout(w[569]));
  fa fa_270 (.a(p[15][22]), .b(p[14][24]), .cin(p[13][26]), .s(w[570]), .cout(w[571]));
  fa fa_271 (.a(p[12][28]), .b(p[11][30]), .cin(p[10][32]), .s(w[572]), .cout(w[573]));
  ha ha_15 (.a(p[9][34]), .b(1'b1), .s(w[574]), .cout(w[575]));
  fa fa_272 (.a(w[575]), .b(w[573]), .cin(w[571]), .s(w[576]), .cout(w[577]));
  fa fa_273 (.a(w[569]), .b(w[567]), .cin(p[16][21]), .s(w[578]), .cout(w[579]));
  fa fa_274 (.a(p[15][23]), .b(p[14][25]), .cin(p[13][27]), .s(w[580]), .cout(w[581]));
  fa fa_275 (.a(p[12][29]), .b(p[11][31]), .cin(p[10][33]), .s(w[582]), .cout(w[583]));
  fa fa_276 (.a(w[583]), .b(w[581]), .cin(w[579]), .s(w[584]), .cout(w[585]));
  fa fa_277 (.a(w[577]), .b(p[16][22]), .cin(p[15][24]), .s(w[586]), .cout(w[587]));
  fa fa_278 (.a(p[14][26]), .b(p[13][28]), .cin(p[12][30]), .s(w[588]), .cout(w[589]));
  fa fa_279 (.a(p[11][32]), .b(p[10][34]), .cin(1'b1), .s(w[590]), .cout(w[591]));
  fa fa_280 (.a(w[591]), .b(w[589]), .cin(w[587]), .s(w[592]), .cout(w[593]));
  fa fa_281 (.a(w[585]), .b(p[16][23]), .cin(p[15][25]), .s(w[594]), .cout(w[595]));
  fa fa_282 (.a(p[14][27]), .b(p[13][29]), .cin(p[12][31]), .s(w[596]), .cout(w[597]));
  ha ha_16 (.a(p[11][33]), .b(p[10][35]), .s(w[598]), .cout(w[599]));
  fa fa_283 (.a(w[599]), .b(w[597]), .cin(w[595]), .s(w[600]), .cout(w[601]));
  fa fa_284 (.a(w[593]), .b(p[16][24]), .cin(p[15][26]), .s(w[602]), .cout(w[603]));
  fa fa_285 (.a(p[14][28]), .b(p[13][30]), .cin(p[12][32]), .s(w[604]), .cout(w[605]));
  ha ha_17 (.a(p[11][34]), .b(1'b1), .s(w[606]), .cout(w[607]));
  fa fa_286 (.a(w[607]), .b(w[605]), .cin(w[603]), .s(w[608]), .cout(w[609]));
  fa fa_287 (.a(w[601]), .b(p[16][25]), .cin(p[15][27]), .s(w[610]), .cout(w[611]));
  fa fa_288 (.a(p[14][29]), .b(p[13][31]), .cin(p[12][33]), .s(w[612]), .cout(w[613]));
  fa fa_289 (.a(w[613]), .b(w[611]), .cin(w[609]), .s(w[614]), .cout(w[615]));
  fa fa_290 (.a(p[16][26]), .b(p[15][28]), .cin(p[14][30]), .s(w[616]), .cout(w[617]));
  fa fa_291 (.a(p[13][32]), .b(p[12][34]), .cin(1'b1), .s(w[618]), .cout(w[619]));
  fa fa_292 (.a(w[619]), .b(w[617]), .cin(w[615]), .s(w[620]), .cout(w[621]));
  fa fa_293 (.a(p[16][27]), .b(p[15][29]), .cin(p[14][31]), .s(w[622]), .cout(w[623]));
  ha ha_18 (.a(p[13][33]), .b(p[12][35]), .s(w[624]), .cout(w[625]));
  fa fa_294 (.a(w[625]), .b(w[623]), .cin(w[621]), .s(w[626]), .cout(w[627]));
  fa fa_295 (.a(p[16][28]), .b(p[15][30]), .cin(p[14][32]), .s(w[628]), .cout(w[629]));
  ha ha_19 (.a(p[13][34]), .b(1'b1), .s(w[630]), .cout(w[631]));
  fa fa_296 (.a(w[631]), .b(w[629]), .cin(w[627]), .s(w[632]), .cout(w[633]));
  fa fa_297 (.a(p[16][29]), .b(p[15][31]), .cin(p[14][33]), .s(w[634]), .cout(w[635]));
  fa fa_298 (.a(w[635]), .b(w[633]), .cin(p[16][30]), .s(w[636]), .cout(w[637]));
  fa fa_299 (.a(p[15][32]), .b(p[14][34]), .cin(1'b1), .s(w[638]), .cout(w[639]));
  fa fa_300 (.a(w[639]), .b(w[637]), .cin(p[16][31]), .s(w[640]), .cout(w[641]));
  ha ha_20 (.a(p[15][33]), .b(p[14][35]), .s(w[642]), .cout(w[643]));
  fa fa_301 (.a(w[643]), .b(w[641]), .cin(p[16][32]), .s(w[644]), .cout(w[645]));
  ha ha_21 (.a(p[15][34]), .b(1'b1), .s(w[646]), .cout(w[647]));
  fa fa_302 (.a(w[647]), .b(w[645]), .cin(p[16][33]), .s(w[648]), .cout(w[649]));
  fa fa_303 (.a(w[649]), .b(p[16][34]), .cin(1'b1), .s(w[650]), .cout(w[651]));
  ha ha_22 (.a(w[651]), .b(p[16][35]), .s(w[652]), .cout(w[653]));
  ha ha_23 (.a(p0[2]), .b(w[4]), .s(w[654]), .cout(w[655]));
  fa fa_304 (.a(w[655]), .b(p0[3]), .cin(w[6]), .s(w[656]), .cout(w[657]));
  fa fa_305 (.a(w[657]), .b(w[10]), .cin(w[8]), .s(w[658]), .cout(w[659]));
  fa fa_306 (.a(w[659]), .b(w[14]), .cin(w[12]), .s(w[660]), .cout(w[661]));
  fa fa_307 (.a(w[661]), .b(p0[6]), .cin(w[18]), .s(w[662]), .cout(w[663]));
  fa fa_308 (.a(w[663]), .b(p0[7]), .cin(w[22]), .s(w[664]), .cout(w[665]));
  fa fa_309 (.a(w[665]), .b(w[28]), .cin(w[26]), .s(w[666]), .cout(w[667]));
  fa fa_310 (.a(w[667]), .b(w[34]), .cin(w[32]), .s(w[668]), .cout(w[669]));
  fa fa_311 (.a(w[669]), .b(p0[10]), .cin(w[40]), .s(w[670]), .cout(w[671]));
  ha ha_24 (.a(w[38]), .b(w[36]), .s(w[672]), .cout(w[673]));
  fa fa_312 (.a(w[673]), .b(w[671]), .cin(p0[11]), .s(w[674]), .cout(w[675]));
  fa fa_313 (.a(w[46]), .b(w[44]), .cin(w[42]), .s(w[676]), .cout(w[677]));
  fa fa_314 (.a(w[677]), .b(w[675]), .cin(w[54]), .s(w[678]), .cout(w[679]));
  fa fa_315 (.a(w[52]), .b(w[50]), .cin(w[48]), .s(w[680]), .cout(w[681]));
  fa fa_316 (.a(w[681]), .b(w[679]), .cin(w[62]), .s(w[682]), .cout(w[683]));
  fa fa_317 (.a(w[60]), .b(w[58]), .cin(w[56]), .s(w[684]), .cout(w[685]));
  fa fa_318 (.a(w[685]), .b(w[683]), .cin(p0[14]), .s(w[686]), .cout(w[687]));
  fa fa_319 (.a(w[70]), .b(w[68]), .cin(w[66]), .s(w[688]), .cout(w[689]));
  fa fa_320 (.a(w[689]), .b(w[687]), .cin(p0[15]), .s(w[690]), .cout(w[691]));
  fa fa_321 (.a(w[78]), .b(w[76]), .cin(w[74]), .s(w[692]), .cout(w[693]));
  fa fa_322 (.a(w[693]), .b(w[691]), .cin(w[88]), .s(w[694]), .cout(w[695]));
  fa fa_323 (.a(w[86]), .b(w[84]), .cin(w[82]), .s(w[696]), .cout(w[697]));
  fa fa_324 (.a(w[697]), .b(w[695]), .cin(w[98]), .s(w[698]), .cout(w[699]));
  fa fa_325 (.a(w[96]), .b(w[94]), .cin(w[92]), .s(w[700]), .cout(w[701]));
  fa fa_326 (.a(w[701]), .b(w[699]), .cin(p0[18]), .s(w[702]), .cout(w[703]));
  fa fa_327 (.a(w[108]), .b(w[106]), .cin(w[104]), .s(w[704]), .cout(w[705]));
  ha ha_25 (.a(w[102]), .b(w[100]), .s(w[706]), .cout(w[707]));
  fa fa_328 (.a(w[707]), .b(w[705]), .cin(w[703]), .s(w[708]), .cout(w[709]));
  fa fa_329 (.a(p0[19]), .b(w[118]), .cin(w[116]), .s(w[710]), .cout(w[711]));
  fa fa_330 (.a(w[114]), .b(w[112]), .cin(w[110]), .s(w[712]), .cout(w[713]));
  fa fa_331 (.a(w[713]), .b(w[711]), .cin(w[709]), .s(w[714]), .cout(w[715]));
  fa fa_332 (.a(w[130]), .b(w[128]), .cin(w[126]), .s(w[716]), .cout(w[717]));
  fa fa_333 (.a(w[124]), .b(w[122]), .cin(w[120]), .s(w[718]), .cout(w[719]));
  fa fa_334 (.a(w[719]), .b(w[717]), .cin(w[715]), .s(w[720]), .cout(w[721]));
  fa fa_335 (.a(w[142]), .b(w[140]), .cin(w[138]), .s(w[722]), .cout(w[723]));
  fa fa_336 (.a(w[136]), .b(w[134]), .cin(w[132]), .s(w[724]), .cout(w[725]));
  fa fa_337 (.a(w[725]), .b(w[723]), .cin(w[721]), .s(w[726]), .cout(w[727]));
  fa fa_338 (.a(p0[22]), .b(w[154]), .cin(w[152]), .s(w[728]), .cout(w[729]));
  fa fa_339 (.a(w[150]), .b(w[148]), .cin(w[146]), .s(w[730]), .cout(w[731]));
  fa fa_340 (.a(w[731]), .b(w[729]), .cin(w[727]), .s(w[732]), .cout(w[733]));
  fa fa_341 (.a(p0[23]), .b(w[166]), .cin(w[164]), .s(w[734]), .cout(w[735]));
  fa fa_342 (.a(w[162]), .b(w[160]), .cin(w[158]), .s(w[736]), .cout(w[737]));
  fa fa_343 (.a(w[737]), .b(w[735]), .cin(w[733]), .s(w[738]), .cout(w[739]));
  fa fa_344 (.a(w[180]), .b(w[178]), .cin(w[176]), .s(w[740]), .cout(w[741]));
  fa fa_345 (.a(w[174]), .b(w[172]), .cin(w[170]), .s(w[742]), .cout(w[743]));
  fa fa_346 (.a(w[743]), .b(w[741]), .cin(w[739]), .s(w[744]), .cout(w[745]));
  fa fa_347 (.a(w[194]), .b(w[192]), .cin(w[190]), .s(w[746]), .cout(w[747]));
  fa fa_348 (.a(w[188]), .b(w[186]), .cin(w[184]), .s(w[748]), .cout(w[749]));
  fa fa_349 (.a(w[749]), .b(w[747]), .cin(w[745]), .s(w[750]), .cout(w[751]));
  fa fa_350 (.a(p0[26]), .b(w[208]), .cin(w[206]), .s(w[752]), .cout(w[753]));
  fa fa_351 (.a(w[204]), .b(w[202]), .cin(w[200]), .s(w[754]), .cout(w[755]));
  ha ha_26 (.a(w[198]), .b(w[196]), .s(w[756]), .cout(w[757]));
  fa fa_352 (.a(w[757]), .b(w[755]), .cin(w[753]), .s(w[758]), .cout(w[759]));
  fa fa_353 (.a(w[751]), .b(p0[27]), .cin(w[222]), .s(w[760]), .cout(w[761]));
  fa fa_354 (.a(w[220]), .b(w[218]), .cin(w[216]), .s(w[762]), .cout(w[763]));
  fa fa_355 (.a(w[214]), .b(w[212]), .cin(w[210]), .s(w[764]), .cout(w[765]));
  fa fa_356 (.a(w[765]), .b(w[763]), .cin(w[761]), .s(w[766]), .cout(w[767]));
  fa fa_357 (.a(w[759]), .b(w[238]), .cin(w[236]), .s(w[768]), .cout(w[769]));
  fa fa_358 (.a(w[234]), .b(w[232]), .cin(w[230]), .s(w[770]), .cout(w[771]));
  fa fa_359 (.a(w[228]), .b(w[226]), .cin(w[224]), .s(w[772]), .cout(w[773]));
  fa fa_360 (.a(w[773]), .b(w[771]), .cin(w[769]), .s(w[774]), .cout(w[775]));
  fa fa_361 (.a(w[767]), .b(w[254]), .cin(w[252]), .s(w[776]), .cout(w[777]));
  fa fa_362 (.a(w[250]), .b(w[248]), .cin(w[246]), .s(w[778]), .cout(w[779]));
  fa fa_363 (.a(w[244]), .b(w[242]), .cin(w[240]), .s(w[780]), .cout(w[781]));
  fa fa_364 (.a(w[781]), .b(w[779]), .cin(w[777]), .s(w[782]), .cout(w[783]));
  fa fa_365 (.a(w[775]), .b(p0[30]), .cin(w[270]), .s(w[784]), .cout(w[785]));
  fa fa_366 (.a(w[268]), .b(w[266]), .cin(w[264]), .s(w[786]), .cout(w[787]));
  fa fa_367 (.a(w[262]), .b(w[260]), .cin(w[258]), .s(w[788]), .cout(w[789]));
  fa fa_368 (.a(w[789]), .b(w[787]), .cin(w[785]), .s(w[790]), .cout(w[791]));
  fa fa_369 (.a(w[783]), .b(p0[31]), .cin(w[286]), .s(w[792]), .cout(w[793]));
  fa fa_370 (.a(w[284]), .b(w[282]), .cin(w[280]), .s(w[794]), .cout(w[795]));
  fa fa_371 (.a(w[278]), .b(w[276]), .cin(w[274]), .s(w[796]), .cout(w[797]));
  fa fa_372 (.a(w[797]), .b(w[795]), .cin(w[793]), .s(w[798]), .cout(w[799]));
  fa fa_373 (.a(w[791]), .b(p0[32]), .cin(w[302]), .s(w[800]), .cout(w[801]));
  fa fa_374 (.a(w[300]), .b(w[298]), .cin(w[296]), .s(w[802]), .cout(w[803]));
  fa fa_375 (.a(w[294]), .b(w[292]), .cin(w[290]), .s(w[804]), .cout(w[805]));
  fa fa_376 (.a(w[805]), .b(w[803]), .cin(w[801]), .s(w[806]), .cout(w[807]));
  fa fa_377 (.a(w[799]), .b(p0[33]), .cin(w[318]), .s(w[808]), .cout(w[809]));
  fa fa_378 (.a(w[316]), .b(w[314]), .cin(w[312]), .s(w[810]), .cout(w[811]));
  fa fa_379 (.a(w[310]), .b(w[308]), .cin(w[306]), .s(w[812]), .cout(w[813]));
  fa fa_380 (.a(w[813]), .b(w[811]), .cin(w[809]), .s(w[814]), .cout(w[815]));
  fa fa_381 (.a(w[807]), .b(p0[34]), .cin(w[334]), .s(w[816]), .cout(w[817]));
  fa fa_382 (.a(w[332]), .b(w[330]), .cin(w[328]), .s(w[818]), .cout(w[819]));
  fa fa_383 (.a(w[326]), .b(w[324]), .cin(w[322]), .s(w[820]), .cout(w[821]));
  fa fa_384 (.a(w[821]), .b(w[819]), .cin(w[817]), .s(w[822]), .cout(w[823]));
  fa fa_385 (.a(w[815]), .b(p0[35]), .cin(w[350]), .s(w[824]), .cout(w[825]));
  fa fa_386 (.a(w[348]), .b(w[346]), .cin(w[344]), .s(w[826]), .cout(w[827]));
  fa fa_387 (.a(w[342]), .b(w[340]), .cin(w[338]), .s(w[828]), .cout(w[829]));
  fa fa_388 (.a(w[829]), .b(w[827]), .cin(w[825]), .s(w[830]), .cout(w[831]));
  fa fa_389 (.a(w[823]), .b(p0[36]), .cin(w[366]), .s(w[832]), .cout(w[833]));
  fa fa_390 (.a(w[364]), .b(w[362]), .cin(w[360]), .s(w[834]), .cout(w[835]));
  fa fa_391 (.a(w[358]), .b(w[356]), .cin(w[354]), .s(w[836]), .cout(w[837]));
  fa fa_392 (.a(w[837]), .b(w[835]), .cin(w[833]), .s(w[838]), .cout(w[839]));
  fa fa_393 (.a(w[831]), .b(p0[37]), .cin(w[382]), .s(w[840]), .cout(w[841]));
  fa fa_394 (.a(w[380]), .b(w[378]), .cin(w[376]), .s(w[842]), .cout(w[843]));
  fa fa_395 (.a(w[374]), .b(w[372]), .cin(w[370]), .s(w[844]), .cout(w[845]));
  fa fa_396 (.a(w[845]), .b(w[843]), .cin(w[841]), .s(w[846]), .cout(w[847]));
  fa fa_397 (.a(w[839]), .b(w[398]), .cin(w[396]), .s(w[848]), .cout(w[849]));
  fa fa_398 (.a(w[394]), .b(w[392]), .cin(w[390]), .s(w[850]), .cout(w[851]));
  fa fa_399 (.a(w[388]), .b(w[386]), .cin(w[384]), .s(w[852]), .cout(w[853]));
  fa fa_400 (.a(w[853]), .b(w[851]), .cin(w[849]), .s(w[854]), .cout(w[855]));
  fa fa_401 (.a(w[847]), .b(w[414]), .cin(w[412]), .s(w[856]), .cout(w[857]));
  fa fa_402 (.a(w[410]), .b(w[408]), .cin(w[406]), .s(w[858]), .cout(w[859]));
  fa fa_403 (.a(w[404]), .b(w[402]), .cin(w[400]), .s(w[860]), .cout(w[861]));
  fa fa_404 (.a(w[861]), .b(w[859]), .cin(w[857]), .s(w[862]), .cout(w[863]));
  fa fa_405 (.a(w[855]), .b(w[430]), .cin(w[428]), .s(w[864]), .cout(w[865]));
  fa fa_406 (.a(w[426]), .b(w[424]), .cin(w[422]), .s(w[866]), .cout(w[867]));
  fa fa_407 (.a(w[420]), .b(w[418]), .cin(w[416]), .s(w[868]), .cout(w[869]));
  fa fa_408 (.a(w[869]), .b(w[867]), .cin(w[865]), .s(w[870]), .cout(w[871]));
  fa fa_409 (.a(w[863]), .b(p[3][35]), .cin(w[444]), .s(w[872]), .cout(w[873]));
  fa fa_410 (.a(w[442]), .b(w[440]), .cin(w[438]), .s(w[874]), .cout(w[875]));
  fa fa_411 (.a(w[436]), .b(w[434]), .cin(w[432]), .s(w[876]), .cout(w[877]));
  fa fa_412 (.a(w[877]), .b(w[875]), .cin(w[873]), .s(w[878]), .cout(w[879]));
  fa fa_413 (.a(w[871]), .b(w[458]), .cin(w[456]), .s(w[880]), .cout(w[881]));
  fa fa_414 (.a(w[454]), .b(w[452]), .cin(w[450]), .s(w[882]), .cout(w[883]));
  ha ha_27 (.a(w[448]), .b(w[446]), .s(w[884]), .cout(w[885]));
  fa fa_415 (.a(w[885]), .b(w[883]), .cin(w[881]), .s(w[886]), .cout(w[887]));
  fa fa_416 (.a(w[879]), .b(w[472]), .cin(w[470]), .s(w[888]), .cout(w[889]));
  fa fa_417 (.a(w[468]), .b(w[466]), .cin(w[464]), .s(w[890]), .cout(w[891]));
  ha ha_28 (.a(w[462]), .b(w[460]), .s(w[892]), .cout(w[893]));
  fa fa_418 (.a(w[893]), .b(w[891]), .cin(w[889]), .s(w[894]), .cout(w[895]));
  fa fa_419 (.a(w[887]), .b(w[486]), .cin(w[484]), .s(w[896]), .cout(w[897]));
  fa fa_420 (.a(w[482]), .b(w[480]), .cin(w[478]), .s(w[898]), .cout(w[899]));
  ha ha_29 (.a(w[476]), .b(w[474]), .s(w[900]), .cout(w[901]));
  fa fa_421 (.a(w[901]), .b(w[899]), .cin(w[897]), .s(w[902]), .cout(w[903]));
  fa fa_422 (.a(w[895]), .b(p[5][35]), .cin(w[498]), .s(w[904]), .cout(w[905]));
  fa fa_423 (.a(w[496]), .b(w[494]), .cin(w[492]), .s(w[906]), .cout(w[907]));
  ha ha_30 (.a(w[490]), .b(w[488]), .s(w[908]), .cout(w[909]));
  fa fa_424 (.a(w[909]), .b(w[907]), .cin(w[905]), .s(w[910]), .cout(w[911]));
  fa fa_425 (.a(w[903]), .b(w[510]), .cin(w[508]), .s(w[912]), .cout(w[913]));
  fa fa_426 (.a(w[506]), .b(w[504]), .cin(w[502]), .s(w[914]), .cout(w[915]));
  fa fa_427 (.a(w[915]), .b(w[913]), .cin(w[911]), .s(w[916]), .cout(w[917]));
  fa fa_428 (.a(w[522]), .b(w[520]), .cin(w[518]), .s(w[918]), .cout(w[919]));
  fa fa_429 (.a(w[516]), .b(w[514]), .cin(w[512]), .s(w[920]), .cout(w[921]));
  fa fa_430 (.a(w[921]), .b(w[919]), .cin(w[917]), .s(w[922]), .cout(w[923]));
  fa fa_431 (.a(w[534]), .b(w[532]), .cin(w[530]), .s(w[924]), .cout(w[925]));
  fa fa_432 (.a(w[528]), .b(w[526]), .cin(w[524]), .s(w[926]), .cout(w[927]));
  fa fa_433 (.a(w[927]), .b(w[925]), .cin(w[923]), .s(w[928]), .cout(w[929]));
  fa fa_434 (.a(p[7][35]), .b(w[544]), .cin(w[542]), .s(w[930]), .cout(w[931]));
  fa fa_435 (.a(w[540]), .b(w[538]), .cin(w[536]), .s(w[932]), .cout(w[933]));
  fa fa_436 (.a(w[933]), .b(w[931]), .cin(w[929]), .s(w[934]), .cout(w[935]));
  fa fa_437 (.a(w[554]), .b(w[552]), .cin(w[550]), .s(w[936]), .cout(w[937]));
  ha ha_31 (.a(w[548]), .b(w[546]), .s(w[938]), .cout(w[939]));
  fa fa_438 (.a(w[939]), .b(w[937]), .cin(w[935]), .s(w[940]), .cout(w[941]));
  fa fa_439 (.a(w[564]), .b(w[562]), .cin(w[560]), .s(w[942]), .cout(w[943]));
  ha ha_32 (.a(w[558]), .b(w[556]), .s(w[944]), .cout(w[945]));
  fa fa_440 (.a(w[945]), .b(w[943]), .cin(w[941]), .s(w[946]), .cout(w[947]));
  fa fa_441 (.a(w[574]), .b(w[572]), .cin(w[570]), .s(w[948]), .cout(w[949]));
  ha ha_33 (.a(w[568]), .b(w[566]), .s(w[950]), .cout(w[951]));
  fa fa_442 (.a(w[951]), .b(w[949]), .cin(w[947]), .s(w[952]), .cout(w[953]));
  fa fa_443 (.a(p[9][35]), .b(w[582]), .cin(w[580]), .s(w[954]), .cout(w[955]));
  ha ha_34 (.a(w[578]), .b(w[576]), .s(w[956]), .cout(w[957]));
  fa fa_444 (.a(w[957]), .b(w[955]), .cin(w[953]), .s(w[958]), .cout(w[959]));
  fa fa_445 (.a(w[590]), .b(w[588]), .cin(w[586]), .s(w[960]), .cout(w[961]));
  fa fa_446 (.a(w[961]), .b(w[959]), .cin(w[598]), .s(w[962]), .cout(w[963]));
  fa fa_447 (.a(w[596]), .b(w[594]), .cin(w[592]), .s(w[964]), .cout(w[965]));
  fa fa_448 (.a(w[965]), .b(w[963]), .cin(w[606]), .s(w[966]), .cout(w[967]));
  fa fa_449 (.a(w[604]), .b(w[602]), .cin(w[600]), .s(w[968]), .cout(w[969]));
  fa fa_450 (.a(w[969]), .b(w[967]), .cin(p[11][35]), .s(w[970]), .cout(w[971]));
  fa fa_451 (.a(w[612]), .b(w[610]), .cin(w[608]), .s(w[972]), .cout(w[973]));
  fa fa_452 (.a(w[973]), .b(w[971]), .cin(w[618]), .s(w[974]), .cout(w[975]));
  ha ha_35 (.a(w[616]), .b(w[614]), .s(w[976]), .cout(w[977]));
  fa fa_453 (.a(w[977]), .b(w[975]), .cin(w[624]), .s(w[978]), .cout(w[979]));
  ha ha_36 (.a(w[622]), .b(w[620]), .s(w[980]), .cout(w[981]));
  fa fa_454 (.a(w[981]), .b(w[979]), .cin(w[630]), .s(w[982]), .cout(w[983]));
  ha ha_37 (.a(w[628]), .b(w[626]), .s(w[984]), .cout(w[985]));
  fa fa_455 (.a(w[985]), .b(w[983]), .cin(p[13][35]), .s(w[986]), .cout(w[987]));
  ha ha_38 (.a(w[634]), .b(w[632]), .s(w[988]), .cout(w[989]));
  fa fa_456 (.a(w[989]), .b(w[987]), .cin(w[638]), .s(w[990]), .cout(w[991]));
  fa fa_457 (.a(w[991]), .b(w[642]), .cin(w[640]), .s(w[992]), .cout(w[993]));
  fa fa_458 (.a(w[993]), .b(w[646]), .cin(w[644]), .s(w[994]), .cout(w[995]));
  fa fa_459 (.a(w[995]), .b(p[15][35]), .cin(w[648]), .s(w[996]), .cout(w[997]));
  ha ha_39 (.a(w[997]), .b(w[650]), .s(w[998]), .cout(w[999]));
  ha ha_40 (.a(w[999]), .b(w[652]), .s(w[1000]), .cout(w[1001]));
  ha ha_41 (.a(w[16]), .b(w[662]), .s(w[1002]), .cout(w[1003]));
  fa fa_460 (.a(w[1003]), .b(w[20]), .cin(w[664]), .s(w[1004]), .cout(w[1005]));
  fa fa_461 (.a(w[1005]), .b(w[24]), .cin(w[666]), .s(w[1006]), .cout(w[1007]));
  fa fa_462 (.a(w[1007]), .b(w[30]), .cin(w[668]), .s(w[1008]), .cout(w[1009]));
  fa fa_463 (.a(w[1009]), .b(w[672]), .cin(w[670]), .s(w[1010]), .cout(w[1011]));
  fa fa_464 (.a(w[1011]), .b(w[676]), .cin(w[674]), .s(w[1012]), .cout(w[1013]));
  fa fa_465 (.a(w[1013]), .b(w[680]), .cin(w[678]), .s(w[1014]), .cout(w[1015]));
  fa fa_466 (.a(w[1015]), .b(w[684]), .cin(w[682]), .s(w[1016]), .cout(w[1017]));
  fa fa_467 (.a(w[1017]), .b(w[64]), .cin(w[688]), .s(w[1018]), .cout(w[1019]));
  fa fa_468 (.a(w[1019]), .b(w[72]), .cin(w[692]), .s(w[1020]), .cout(w[1021]));
  fa fa_469 (.a(w[1021]), .b(w[80]), .cin(w[696]), .s(w[1022]), .cout(w[1023]));
  fa fa_470 (.a(w[1023]), .b(w[90]), .cin(w[700]), .s(w[1024]), .cout(w[1025]));
  fa fa_471 (.a(w[1025]), .b(w[706]), .cin(w[704]), .s(w[1026]), .cout(w[1027]));
  fa fa_472 (.a(w[1027]), .b(w[712]), .cin(w[710]), .s(w[1028]), .cout(w[1029]));
  fa fa_473 (.a(w[1029]), .b(w[718]), .cin(w[716]), .s(w[1030]), .cout(w[1031]));
  fa fa_474 (.a(w[1031]), .b(w[724]), .cin(w[722]), .s(w[1032]), .cout(w[1033]));
  fa fa_475 (.a(w[1033]), .b(w[144]), .cin(w[730]), .s(w[1034]), .cout(w[1035]));
  ha ha_42 (.a(w[728]), .b(w[726]), .s(w[1036]), .cout(w[1037]));
  fa fa_476 (.a(w[1037]), .b(w[1035]), .cin(w[156]), .s(w[1038]), .cout(w[1039]));
  fa fa_477 (.a(w[736]), .b(w[734]), .cin(w[732]), .s(w[1040]), .cout(w[1041]));
  fa fa_478 (.a(w[1041]), .b(w[1039]), .cin(w[168]), .s(w[1042]), .cout(w[1043]));
  fa fa_479 (.a(w[742]), .b(w[740]), .cin(w[738]), .s(w[1044]), .cout(w[1045]));
  fa fa_480 (.a(w[1045]), .b(w[1043]), .cin(w[182]), .s(w[1046]), .cout(w[1047]));
  fa fa_481 (.a(w[748]), .b(w[746]), .cin(w[744]), .s(w[1048]), .cout(w[1049]));
  fa fa_482 (.a(w[1049]), .b(w[1047]), .cin(w[756]), .s(w[1050]), .cout(w[1051]));
  fa fa_483 (.a(w[754]), .b(w[752]), .cin(w[750]), .s(w[1052]), .cout(w[1053]));
  fa fa_484 (.a(w[1053]), .b(w[1051]), .cin(w[764]), .s(w[1054]), .cout(w[1055]));
  fa fa_485 (.a(w[762]), .b(w[760]), .cin(w[758]), .s(w[1056]), .cout(w[1057]));
  fa fa_486 (.a(w[1057]), .b(w[1055]), .cin(w[772]), .s(w[1058]), .cout(w[1059]));
  fa fa_487 (.a(w[770]), .b(w[768]), .cin(w[766]), .s(w[1060]), .cout(w[1061]));
  fa fa_488 (.a(w[1061]), .b(w[1059]), .cin(w[780]), .s(w[1062]), .cout(w[1063]));
  fa fa_489 (.a(w[778]), .b(w[776]), .cin(w[774]), .s(w[1064]), .cout(w[1065]));
  fa fa_490 (.a(w[1065]), .b(w[1063]), .cin(w[256]), .s(w[1066]), .cout(w[1067]));
  fa fa_491 (.a(w[788]), .b(w[786]), .cin(w[784]), .s(w[1068]), .cout(w[1069]));
  fa fa_492 (.a(w[1069]), .b(w[1067]), .cin(w[272]), .s(w[1070]), .cout(w[1071]));
  fa fa_493 (.a(w[796]), .b(w[794]), .cin(w[792]), .s(w[1072]), .cout(w[1073]));
  fa fa_494 (.a(w[1073]), .b(w[1071]), .cin(w[288]), .s(w[1074]), .cout(w[1075]));
  fa fa_495 (.a(w[804]), .b(w[802]), .cin(w[800]), .s(w[1076]), .cout(w[1077]));
  fa fa_496 (.a(w[1077]), .b(w[1075]), .cin(w[304]), .s(w[1078]), .cout(w[1079]));
  fa fa_497 (.a(w[812]), .b(w[810]), .cin(w[808]), .s(w[1080]), .cout(w[1081]));
  fa fa_498 (.a(w[1081]), .b(w[1079]), .cin(w[320]), .s(w[1082]), .cout(w[1083]));
  fa fa_499 (.a(w[820]), .b(w[818]), .cin(w[816]), .s(w[1084]), .cout(w[1085]));
  fa fa_500 (.a(w[1085]), .b(w[1083]), .cin(w[336]), .s(w[1086]), .cout(w[1087]));
  fa fa_501 (.a(w[828]), .b(w[826]), .cin(w[824]), .s(w[1088]), .cout(w[1089]));
  fa fa_502 (.a(w[1089]), .b(w[1087]), .cin(w[352]), .s(w[1090]), .cout(w[1091]));
  fa fa_503 (.a(w[836]), .b(w[834]), .cin(w[832]), .s(w[1092]), .cout(w[1093]));
  fa fa_504 (.a(w[1093]), .b(w[1091]), .cin(w[368]), .s(w[1094]), .cout(w[1095]));
  fa fa_505 (.a(w[844]), .b(w[842]), .cin(w[840]), .s(w[1096]), .cout(w[1097]));
  fa fa_506 (.a(w[1097]), .b(w[1095]), .cin(w[852]), .s(w[1098]), .cout(w[1099]));
  fa fa_507 (.a(w[850]), .b(w[848]), .cin(w[846]), .s(w[1100]), .cout(w[1101]));
  fa fa_508 (.a(w[1101]), .b(w[1099]), .cin(w[860]), .s(w[1102]), .cout(w[1103]));
  fa fa_509 (.a(w[858]), .b(w[856]), .cin(w[854]), .s(w[1104]), .cout(w[1105]));
  fa fa_510 (.a(w[1105]), .b(w[1103]), .cin(w[868]), .s(w[1106]), .cout(w[1107]));
  fa fa_511 (.a(w[866]), .b(w[864]), .cin(w[862]), .s(w[1108]), .cout(w[1109]));
  fa fa_512 (.a(w[1109]), .b(w[1107]), .cin(w[876]), .s(w[1110]), .cout(w[1111]));
  fa fa_513 (.a(w[874]), .b(w[872]), .cin(w[870]), .s(w[1112]), .cout(w[1113]));
  fa fa_514 (.a(w[1113]), .b(w[1111]), .cin(w[884]), .s(w[1114]), .cout(w[1115]));
  fa fa_515 (.a(w[882]), .b(w[880]), .cin(w[878]), .s(w[1116]), .cout(w[1117]));
  fa fa_516 (.a(w[1117]), .b(w[1115]), .cin(w[892]), .s(w[1118]), .cout(w[1119]));
  fa fa_517 (.a(w[890]), .b(w[888]), .cin(w[886]), .s(w[1120]), .cout(w[1121]));
  fa fa_518 (.a(w[1121]), .b(w[1119]), .cin(w[900]), .s(w[1122]), .cout(w[1123]));
  fa fa_519 (.a(w[898]), .b(w[896]), .cin(w[894]), .s(w[1124]), .cout(w[1125]));
  fa fa_520 (.a(w[1125]), .b(w[1123]), .cin(w[908]), .s(w[1126]), .cout(w[1127]));
  fa fa_521 (.a(w[906]), .b(w[904]), .cin(w[902]), .s(w[1128]), .cout(w[1129]));
  fa fa_522 (.a(w[1129]), .b(w[1127]), .cin(w[500]), .s(w[1130]), .cout(w[1131]));
  fa fa_523 (.a(w[914]), .b(w[912]), .cin(w[910]), .s(w[1132]), .cout(w[1133]));
  fa fa_524 (.a(w[1133]), .b(w[1131]), .cin(w[920]), .s(w[1134]), .cout(w[1135]));
  ha ha_43 (.a(w[918]), .b(w[916]), .s(w[1136]), .cout(w[1137]));
  fa fa_525 (.a(w[1137]), .b(w[1135]), .cin(w[926]), .s(w[1138]), .cout(w[1139]));
  ha ha_44 (.a(w[924]), .b(w[922]), .s(w[1140]), .cout(w[1141]));
  fa fa_526 (.a(w[1141]), .b(w[1139]), .cin(w[932]), .s(w[1142]), .cout(w[1143]));
  ha ha_45 (.a(w[930]), .b(w[928]), .s(w[1144]), .cout(w[1145]));
  fa fa_527 (.a(w[1145]), .b(w[1143]), .cin(w[938]), .s(w[1146]), .cout(w[1147]));
  ha ha_46 (.a(w[936]), .b(w[934]), .s(w[1148]), .cout(w[1149]));
  fa fa_528 (.a(w[1149]), .b(w[1147]), .cin(w[944]), .s(w[1150]), .cout(w[1151]));
  ha ha_47 (.a(w[942]), .b(w[940]), .s(w[1152]), .cout(w[1153]));
  fa fa_529 (.a(w[1153]), .b(w[1151]), .cin(w[950]), .s(w[1154]), .cout(w[1155]));
  ha ha_48 (.a(w[948]), .b(w[946]), .s(w[1156]), .cout(w[1157]));
  fa fa_530 (.a(w[1157]), .b(w[1155]), .cin(w[956]), .s(w[1158]), .cout(w[1159]));
  ha ha_49 (.a(w[954]), .b(w[952]), .s(w[1160]), .cout(w[1161]));
  fa fa_531 (.a(w[1161]), .b(w[1159]), .cin(w[584]), .s(w[1162]), .cout(w[1163]));
  ha ha_50 (.a(w[960]), .b(w[958]), .s(w[1164]), .cout(w[1165]));
  fa fa_532 (.a(w[1165]), .b(w[1163]), .cin(w[964]), .s(w[1166]), .cout(w[1167]));
  fa fa_533 (.a(w[1167]), .b(w[968]), .cin(w[966]), .s(w[1168]), .cout(w[1169]));
  fa fa_534 (.a(w[1169]), .b(w[972]), .cin(w[970]), .s(w[1170]), .cout(w[1171]));
  fa fa_535 (.a(w[1171]), .b(w[976]), .cin(w[974]), .s(w[1172]), .cout(w[1173]));
  fa fa_536 (.a(w[1173]), .b(w[980]), .cin(w[978]), .s(w[1174]), .cout(w[1175]));
  fa fa_537 (.a(w[1175]), .b(w[984]), .cin(w[982]), .s(w[1176]), .cout(w[1177]));
  fa fa_538 (.a(w[1177]), .b(w[988]), .cin(w[986]), .s(w[1178]), .cout(w[1179]));
  fa fa_539 (.a(w[1179]), .b(w[636]), .cin(w[990]), .s(w[1180]), .cout(w[1181]));
  ha ha_51 (.a(w[1181]), .b(w[992]), .s(w[1182]), .cout(w[1183]));
  ha ha_52 (.a(w[1183]), .b(w[994]), .s(w[1184]), .cout(w[1185]));
  ha ha_53 (.a(w[1185]), .b(w[996]), .s(w[1186]), .cout(w[1187]));
  ha ha_54 (.a(w[1187]), .b(w[998]), .s(w[1188]), .cout(w[1189]));
  ha ha_55 (.a(w[1189]), .b(w[1000]), .s(w[1190]), .cout(w[1191]));
  ha ha_56 (.a(w[686]), .b(w[1018]), .s(w[1192]), .cout(w[1193]));
  fa fa_540 (.a(w[1193]), .b(w[690]), .cin(w[1020]), .s(w[1194]), .cout(w[1195]));
  fa fa_541 (.a(w[1195]), .b(w[694]), .cin(w[1022]), .s(w[1196]), .cout(w[1197]));
  fa fa_542 (.a(w[1197]), .b(w[698]), .cin(w[1024]), .s(w[1198]), .cout(w[1199]));
  fa fa_543 (.a(w[1199]), .b(w[702]), .cin(w[1026]), .s(w[1200]), .cout(w[1201]));
  fa fa_544 (.a(w[1201]), .b(w[708]), .cin(w[1028]), .s(w[1202]), .cout(w[1203]));
  fa fa_545 (.a(w[1203]), .b(w[714]), .cin(w[1030]), .s(w[1204]), .cout(w[1205]));
  fa fa_546 (.a(w[1205]), .b(w[720]), .cin(w[1032]), .s(w[1206]), .cout(w[1207]));
  fa fa_547 (.a(w[1207]), .b(w[1036]), .cin(w[1034]), .s(w[1208]), .cout(w[1209]));
  fa fa_548 (.a(w[1209]), .b(w[1040]), .cin(w[1038]), .s(w[1210]), .cout(w[1211]));
  fa fa_549 (.a(w[1211]), .b(w[1044]), .cin(w[1042]), .s(w[1212]), .cout(w[1213]));
  fa fa_550 (.a(w[1213]), .b(w[1048]), .cin(w[1046]), .s(w[1214]), .cout(w[1215]));
  fa fa_551 (.a(w[1215]), .b(w[1052]), .cin(w[1050]), .s(w[1216]), .cout(w[1217]));
  fa fa_552 (.a(w[1217]), .b(w[1056]), .cin(w[1054]), .s(w[1218]), .cout(w[1219]));
  fa fa_553 (.a(w[1219]), .b(w[1060]), .cin(w[1058]), .s(w[1220]), .cout(w[1221]));
  fa fa_554 (.a(w[1221]), .b(w[1064]), .cin(w[1062]), .s(w[1222]), .cout(w[1223]));
  fa fa_555 (.a(w[1223]), .b(w[782]), .cin(w[1068]), .s(w[1224]), .cout(w[1225]));
  fa fa_556 (.a(w[1225]), .b(w[790]), .cin(w[1072]), .s(w[1226]), .cout(w[1227]));
  fa fa_557 (.a(w[1227]), .b(w[798]), .cin(w[1076]), .s(w[1228]), .cout(w[1229]));
  fa fa_558 (.a(w[1229]), .b(w[806]), .cin(w[1080]), .s(w[1230]), .cout(w[1231]));
  fa fa_559 (.a(w[1231]), .b(w[814]), .cin(w[1084]), .s(w[1232]), .cout(w[1233]));
  fa fa_560 (.a(w[1233]), .b(w[822]), .cin(w[1088]), .s(w[1234]), .cout(w[1235]));
  fa fa_561 (.a(w[1235]), .b(w[830]), .cin(w[1092]), .s(w[1236]), .cout(w[1237]));
  fa fa_562 (.a(w[1237]), .b(w[838]), .cin(w[1096]), .s(w[1238]), .cout(w[1239]));
  fa fa_563 (.a(w[1239]), .b(w[1100]), .cin(w[1098]), .s(w[1240]), .cout(w[1241]));
  fa fa_564 (.a(w[1241]), .b(w[1104]), .cin(w[1102]), .s(w[1242]), .cout(w[1243]));
  fa fa_565 (.a(w[1243]), .b(w[1108]), .cin(w[1106]), .s(w[1244]), .cout(w[1245]));
  fa fa_566 (.a(w[1245]), .b(w[1112]), .cin(w[1110]), .s(w[1246]), .cout(w[1247]));
  fa fa_567 (.a(w[1247]), .b(w[1116]), .cin(w[1114]), .s(w[1248]), .cout(w[1249]));
  fa fa_568 (.a(w[1249]), .b(w[1120]), .cin(w[1118]), .s(w[1250]), .cout(w[1251]));
  fa fa_569 (.a(w[1251]), .b(w[1124]), .cin(w[1122]), .s(w[1252]), .cout(w[1253]));
  fa fa_570 (.a(w[1253]), .b(w[1128]), .cin(w[1126]), .s(w[1254]), .cout(w[1255]));
  fa fa_571 (.a(w[1255]), .b(w[1132]), .cin(w[1130]), .s(w[1256]), .cout(w[1257]));
  fa fa_572 (.a(w[1257]), .b(w[1136]), .cin(w[1134]), .s(w[1258]), .cout(w[1259]));
  fa fa_573 (.a(w[1259]), .b(w[1140]), .cin(w[1138]), .s(w[1260]), .cout(w[1261]));
  fa fa_574 (.a(w[1261]), .b(w[1144]), .cin(w[1142]), .s(w[1262]), .cout(w[1263]));
  fa fa_575 (.a(w[1263]), .b(w[1148]), .cin(w[1146]), .s(w[1264]), .cout(w[1265]));
  fa fa_576 (.a(w[1265]), .b(w[1152]), .cin(w[1150]), .s(w[1266]), .cout(w[1267]));
  fa fa_577 (.a(w[1267]), .b(w[1156]), .cin(w[1154]), .s(w[1268]), .cout(w[1269]));
  fa fa_578 (.a(w[1269]), .b(w[1160]), .cin(w[1158]), .s(w[1270]), .cout(w[1271]));
  fa fa_579 (.a(w[1271]), .b(w[1164]), .cin(w[1162]), .s(w[1272]), .cout(w[1273]));
  fa fa_580 (.a(w[1273]), .b(w[962]), .cin(w[1166]), .s(w[1274]), .cout(w[1275]));
  ha ha_57 (.a(w[1275]), .b(w[1168]), .s(w[1276]), .cout(w[1277]));
  ha ha_58 (.a(w[1277]), .b(w[1170]), .s(w[1278]), .cout(w[1279]));
  ha ha_59 (.a(w[1279]), .b(w[1172]), .s(w[1280]), .cout(w[1281]));
  ha ha_60 (.a(w[1281]), .b(w[1174]), .s(w[1282]), .cout(w[1283]));
  ha ha_61 (.a(w[1283]), .b(w[1176]), .s(w[1284]), .cout(w[1285]));
  ha ha_62 (.a(w[1285]), .b(w[1178]), .s(w[1286]), .cout(w[1287]));
  ha ha_63 (.a(w[1287]), .b(w[1180]), .s(w[1288]), .cout(w[1289]));
  ha ha_64 (.a(w[1289]), .b(w[1182]), .s(w[1290]), .cout(w[1291]));
  ha ha_65 (.a(w[1291]), .b(w[1184]), .s(w[1292]), .cout(w[1293]));
  ha ha_66 (.a(w[1293]), .b(w[1186]), .s(w[1294]), .cout(w[1295]));
  ha ha_67 (.a(w[1295]), .b(w[1188]), .s(w[1296]), .cout(w[1297]));
  ha ha_68 (.a(w[1297]), .b(w[1190]), .s(w[1298]), .cout(w[1299]));
  wire w[1300];
  wire [67:0] row_0 = {w[1298], w[1296], w[1294], w[1292], w[1290], w[1288], w[1286], w[1284], w[1282], w[1280], w[1278], w[1276], w[1274], w[1272], w[1270], w[1268], w[1266], w[1264], w[1262], w[1260], w[1258], w[1256], w[1254], w[1252], w[1250], w[1248], w[1246], w[1244], w[1242], w[1240], w[1094], w[1090], w[1086], w[1082], w[1078], w[1074], w[1070], w[1066], w[1222], w[1220], w[1218], w[1216], w[1214], w[1212], w[1210], w[1208], w[1206], w[1204], w[1202], w[1200], w[1198], w[1196], w[1194], w[1192], w[1016], w[1014], w[1012], w[1010], w[1008], w[1006], w[1004], w[1002], w[660], w[658], w[656], w[654], w[2], w[0]};
  wire [67:0] row_1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, w[1238], w[1236], w[1234], w[1232], w[1230], w[1228], w[1226], w[1224], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
  wire [67:0] prod = row_0 + row_1;

  assign out_prod = prod[63:0];
  assign in_ready = 1;
  assign out_valid = in_valid & ~flush;
endmodule

module fa (
  input a, b, cin,
  output s, cout
);
  assign s = a ^ b ^ cin;
  assign cout = (a & b) | (b & cin) | (a & cin);
endmodule

module ha (
  input a, b,
  output s, cout
);
  assign s = a ^ b;
  assign cout = a & b;
endmodule
